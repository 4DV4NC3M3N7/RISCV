
	
	module Top_module_SV(in,out,sel);
//------------------------------------
//testing functional
			input [31:0]in;
			input [4:0]sel;
			output out;
//------------------------------------

				 ALU();
				 //Register_file();
				 //Data_Memory();
	endmodule
	//*/
	